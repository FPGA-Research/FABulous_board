module template ();
wire Tile_X0Y1_A_I, Tile_X0Y1_A_T, Tile_X0Y1_A_O, Tile_X0Y1_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y1_A (.O(Tile_X0Y1_A_O), .Q(Tile_X0Y1_A_Q), .I(Tile_X0Y1_A_I));

wire Tile_X0Y1_B_I, Tile_X0Y1_B_T, Tile_X0Y1_B_O, Tile_X0Y1_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y1_B (.O(Tile_X0Y1_B_O), .Q(Tile_X0Y1_B_Q), .I(Tile_X0Y1_B_I));

wire Tile_X9Y1_RAM2FAB_D0_O0, Tile_X9Y1_RAM2FAB_D0_O1, Tile_X9Y1_RAM2FAB_D0_O2, Tile_X9Y1_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y1_A (.O0(Tile_X9Y1_RAM2FAB_D0_O0), .O1(Tile_X9Y1_RAM2FAB_D0_O1), .O2(Tile_X9Y1_RAM2FAB_D0_O2), .O3(Tile_X9Y1_RAM2FAB_D0_O3));

wire Tile_X9Y1_RAM2FAB_D1_O0, Tile_X9Y1_RAM2FAB_D1_O1, Tile_X9Y1_RAM2FAB_D1_O2, Tile_X9Y1_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y1_B (.O0(Tile_X9Y1_RAM2FAB_D1_O0), .O1(Tile_X9Y1_RAM2FAB_D1_O1), .O2(Tile_X9Y1_RAM2FAB_D1_O2), .O3(Tile_X9Y1_RAM2FAB_D1_O3));

wire Tile_X9Y1_RAM2FAB_D2_O0, Tile_X9Y1_RAM2FAB_D2_O1, Tile_X9Y1_RAM2FAB_D2_O2, Tile_X9Y1_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y1_C (.O0(Tile_X9Y1_RAM2FAB_D2_O0), .O1(Tile_X9Y1_RAM2FAB_D2_O1), .O2(Tile_X9Y1_RAM2FAB_D2_O2), .O3(Tile_X9Y1_RAM2FAB_D2_O3));

wire Tile_X9Y1_RAM2FAB_D3_O0, Tile_X9Y1_RAM2FAB_D3_O1, Tile_X9Y1_RAM2FAB_D3_O2, Tile_X9Y1_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y1_D (.O0(Tile_X9Y1_RAM2FAB_D3_O0), .O1(Tile_X9Y1_RAM2FAB_D3_O1), .O2(Tile_X9Y1_RAM2FAB_D3_O2), .O3(Tile_X9Y1_RAM2FAB_D3_O3));

wire Tile_X9Y1_FAB2RAM_D0_I0, Tile_X9Y1_FAB2RAM_D0_I1, Tile_X9Y1_FAB2RAM_D0_I2, Tile_X9Y1_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_E (.I0(Tile_X9Y1_FAB2RAM_D0_I0), .I1(Tile_X9Y1_FAB2RAM_D0_I1), .I2(Tile_X9Y1_FAB2RAM_D0_I2), .I3(Tile_X9Y1_FAB2RAM_D0_I3));

wire Tile_X9Y1_FAB2RAM_D1_I0, Tile_X9Y1_FAB2RAM_D1_I1, Tile_X9Y1_FAB2RAM_D1_I2, Tile_X9Y1_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_F (.I0(Tile_X9Y1_FAB2RAM_D1_I0), .I1(Tile_X9Y1_FAB2RAM_D1_I1), .I2(Tile_X9Y1_FAB2RAM_D1_I2), .I3(Tile_X9Y1_FAB2RAM_D1_I3));

wire Tile_X9Y1_FAB2RAM_D2_I0, Tile_X9Y1_FAB2RAM_D2_I1, Tile_X9Y1_FAB2RAM_D2_I2, Tile_X9Y1_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_G (.I0(Tile_X9Y1_FAB2RAM_D2_I0), .I1(Tile_X9Y1_FAB2RAM_D2_I1), .I2(Tile_X9Y1_FAB2RAM_D2_I2), .I3(Tile_X9Y1_FAB2RAM_D2_I3));

wire Tile_X9Y1_FAB2RAM_D3_I0, Tile_X9Y1_FAB2RAM_D3_I1, Tile_X9Y1_FAB2RAM_D3_I2, Tile_X9Y1_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_H (.I0(Tile_X9Y1_FAB2RAM_D3_I0), .I1(Tile_X9Y1_FAB2RAM_D3_I1), .I2(Tile_X9Y1_FAB2RAM_D3_I2), .I3(Tile_X9Y1_FAB2RAM_D3_I3));

wire Tile_X9Y1_FAB2RAM_A0_I0, Tile_X9Y1_FAB2RAM_A0_I1, Tile_X9Y1_FAB2RAM_A0_I2, Tile_X9Y1_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_I (.I0(Tile_X9Y1_FAB2RAM_A0_I0), .I1(Tile_X9Y1_FAB2RAM_A0_I1), .I2(Tile_X9Y1_FAB2RAM_A0_I2), .I3(Tile_X9Y1_FAB2RAM_A0_I3));

wire Tile_X9Y1_FAB2RAM_A1_I0, Tile_X9Y1_FAB2RAM_A1_I1, Tile_X9Y1_FAB2RAM_A1_I2, Tile_X9Y1_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_J (.I0(Tile_X9Y1_FAB2RAM_A1_I0), .I1(Tile_X9Y1_FAB2RAM_A1_I1), .I2(Tile_X9Y1_FAB2RAM_A1_I2), .I3(Tile_X9Y1_FAB2RAM_A1_I3));

wire Tile_X9Y1_FAB2RAM_C_I0, Tile_X9Y1_FAB2RAM_C_I1, Tile_X9Y1_FAB2RAM_C_I2, Tile_X9Y1_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_K (.I0(Tile_X9Y1_FAB2RAM_C_I0), .I1(Tile_X9Y1_FAB2RAM_C_I1), .I2(Tile_X9Y1_FAB2RAM_C_I2), .I3(Tile_X9Y1_FAB2RAM_C_I3));

wire Tile_X0Y2_A_I, Tile_X0Y2_A_T, Tile_X0Y2_A_O, Tile_X0Y2_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y2_A (.O(Tile_X0Y2_A_O), .Q(Tile_X0Y2_A_Q), .I(Tile_X0Y2_A_I));

wire Tile_X0Y2_B_I, Tile_X0Y2_B_T, Tile_X0Y2_B_O, Tile_X0Y2_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y2_B (.O(Tile_X0Y2_B_O), .Q(Tile_X0Y2_B_Q), .I(Tile_X0Y2_B_I));

wire Tile_X9Y2_RAM2FAB_D0_O0, Tile_X9Y2_RAM2FAB_D0_O1, Tile_X9Y2_RAM2FAB_D0_O2, Tile_X9Y2_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y2_A (.O0(Tile_X9Y2_RAM2FAB_D0_O0), .O1(Tile_X9Y2_RAM2FAB_D0_O1), .O2(Tile_X9Y2_RAM2FAB_D0_O2), .O3(Tile_X9Y2_RAM2FAB_D0_O3));

wire Tile_X9Y2_RAM2FAB_D1_O0, Tile_X9Y2_RAM2FAB_D1_O1, Tile_X9Y2_RAM2FAB_D1_O2, Tile_X9Y2_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y2_B (.O0(Tile_X9Y2_RAM2FAB_D1_O0), .O1(Tile_X9Y2_RAM2FAB_D1_O1), .O2(Tile_X9Y2_RAM2FAB_D1_O2), .O3(Tile_X9Y2_RAM2FAB_D1_O3));

wire Tile_X9Y2_RAM2FAB_D2_O0, Tile_X9Y2_RAM2FAB_D2_O1, Tile_X9Y2_RAM2FAB_D2_O2, Tile_X9Y2_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y2_C (.O0(Tile_X9Y2_RAM2FAB_D2_O0), .O1(Tile_X9Y2_RAM2FAB_D2_O1), .O2(Tile_X9Y2_RAM2FAB_D2_O2), .O3(Tile_X9Y2_RAM2FAB_D2_O3));

wire Tile_X9Y2_RAM2FAB_D3_O0, Tile_X9Y2_RAM2FAB_D3_O1, Tile_X9Y2_RAM2FAB_D3_O2, Tile_X9Y2_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y2_D (.O0(Tile_X9Y2_RAM2FAB_D3_O0), .O1(Tile_X9Y2_RAM2FAB_D3_O1), .O2(Tile_X9Y2_RAM2FAB_D3_O2), .O3(Tile_X9Y2_RAM2FAB_D3_O3));

wire Tile_X9Y2_FAB2RAM_D0_I0, Tile_X9Y2_FAB2RAM_D0_I1, Tile_X9Y2_FAB2RAM_D0_I2, Tile_X9Y2_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_E (.I0(Tile_X9Y2_FAB2RAM_D0_I0), .I1(Tile_X9Y2_FAB2RAM_D0_I1), .I2(Tile_X9Y2_FAB2RAM_D0_I2), .I3(Tile_X9Y2_FAB2RAM_D0_I3));

wire Tile_X9Y2_FAB2RAM_D1_I0, Tile_X9Y2_FAB2RAM_D1_I1, Tile_X9Y2_FAB2RAM_D1_I2, Tile_X9Y2_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_F (.I0(Tile_X9Y2_FAB2RAM_D1_I0), .I1(Tile_X9Y2_FAB2RAM_D1_I1), .I2(Tile_X9Y2_FAB2RAM_D1_I2), .I3(Tile_X9Y2_FAB2RAM_D1_I3));

wire Tile_X9Y2_FAB2RAM_D2_I0, Tile_X9Y2_FAB2RAM_D2_I1, Tile_X9Y2_FAB2RAM_D2_I2, Tile_X9Y2_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_G (.I0(Tile_X9Y2_FAB2RAM_D2_I0), .I1(Tile_X9Y2_FAB2RAM_D2_I1), .I2(Tile_X9Y2_FAB2RAM_D2_I2), .I3(Tile_X9Y2_FAB2RAM_D2_I3));

wire Tile_X9Y2_FAB2RAM_D3_I0, Tile_X9Y2_FAB2RAM_D3_I1, Tile_X9Y2_FAB2RAM_D3_I2, Tile_X9Y2_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_H (.I0(Tile_X9Y2_FAB2RAM_D3_I0), .I1(Tile_X9Y2_FAB2RAM_D3_I1), .I2(Tile_X9Y2_FAB2RAM_D3_I2), .I3(Tile_X9Y2_FAB2RAM_D3_I3));

wire Tile_X9Y2_FAB2RAM_A0_I0, Tile_X9Y2_FAB2RAM_A0_I1, Tile_X9Y2_FAB2RAM_A0_I2, Tile_X9Y2_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_I (.I0(Tile_X9Y2_FAB2RAM_A0_I0), .I1(Tile_X9Y2_FAB2RAM_A0_I1), .I2(Tile_X9Y2_FAB2RAM_A0_I2), .I3(Tile_X9Y2_FAB2RAM_A0_I3));

wire Tile_X9Y2_FAB2RAM_A1_I0, Tile_X9Y2_FAB2RAM_A1_I1, Tile_X9Y2_FAB2RAM_A1_I2, Tile_X9Y2_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_J (.I0(Tile_X9Y2_FAB2RAM_A1_I0), .I1(Tile_X9Y2_FAB2RAM_A1_I1), .I2(Tile_X9Y2_FAB2RAM_A1_I2), .I3(Tile_X9Y2_FAB2RAM_A1_I3));

wire Tile_X9Y2_FAB2RAM_C_I0, Tile_X9Y2_FAB2RAM_C_I1, Tile_X9Y2_FAB2RAM_C_I2, Tile_X9Y2_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y2_K (.I0(Tile_X9Y2_FAB2RAM_C_I0), .I1(Tile_X9Y2_FAB2RAM_C_I1), .I2(Tile_X9Y2_FAB2RAM_C_I2), .I3(Tile_X9Y2_FAB2RAM_C_I3));

wire Tile_X0Y3_A_I, Tile_X0Y3_A_T, Tile_X0Y3_A_O, Tile_X0Y3_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y3_A (.O(Tile_X0Y3_A_O), .Q(Tile_X0Y3_A_Q), .I(Tile_X0Y3_A_I));

wire Tile_X0Y3_B_I, Tile_X0Y3_B_T, Tile_X0Y3_B_O, Tile_X0Y3_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y3_B (.O(Tile_X0Y3_B_O), .Q(Tile_X0Y3_B_Q), .I(Tile_X0Y3_B_I));

wire Tile_X9Y3_RAM2FAB_D0_O0, Tile_X9Y3_RAM2FAB_D0_O1, Tile_X9Y3_RAM2FAB_D0_O2, Tile_X9Y3_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y3_A (.O0(Tile_X9Y3_RAM2FAB_D0_O0), .O1(Tile_X9Y3_RAM2FAB_D0_O1), .O2(Tile_X9Y3_RAM2FAB_D0_O2), .O3(Tile_X9Y3_RAM2FAB_D0_O3));

wire Tile_X9Y3_RAM2FAB_D1_O0, Tile_X9Y3_RAM2FAB_D1_O1, Tile_X9Y3_RAM2FAB_D1_O2, Tile_X9Y3_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y3_B (.O0(Tile_X9Y3_RAM2FAB_D1_O0), .O1(Tile_X9Y3_RAM2FAB_D1_O1), .O2(Tile_X9Y3_RAM2FAB_D1_O2), .O3(Tile_X9Y3_RAM2FAB_D1_O3));

wire Tile_X9Y3_RAM2FAB_D2_O0, Tile_X9Y3_RAM2FAB_D2_O1, Tile_X9Y3_RAM2FAB_D2_O2, Tile_X9Y3_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y3_C (.O0(Tile_X9Y3_RAM2FAB_D2_O0), .O1(Tile_X9Y3_RAM2FAB_D2_O1), .O2(Tile_X9Y3_RAM2FAB_D2_O2), .O3(Tile_X9Y3_RAM2FAB_D2_O3));

wire Tile_X9Y3_RAM2FAB_D3_O0, Tile_X9Y3_RAM2FAB_D3_O1, Tile_X9Y3_RAM2FAB_D3_O2, Tile_X9Y3_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y3_D (.O0(Tile_X9Y3_RAM2FAB_D3_O0), .O1(Tile_X9Y3_RAM2FAB_D3_O1), .O2(Tile_X9Y3_RAM2FAB_D3_O2), .O3(Tile_X9Y3_RAM2FAB_D3_O3));

wire Tile_X9Y3_FAB2RAM_D0_I0, Tile_X9Y3_FAB2RAM_D0_I1, Tile_X9Y3_FAB2RAM_D0_I2, Tile_X9Y3_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_E (.I0(Tile_X9Y3_FAB2RAM_D0_I0), .I1(Tile_X9Y3_FAB2RAM_D0_I1), .I2(Tile_X9Y3_FAB2RAM_D0_I2), .I3(Tile_X9Y3_FAB2RAM_D0_I3));

wire Tile_X9Y3_FAB2RAM_D1_I0, Tile_X9Y3_FAB2RAM_D1_I1, Tile_X9Y3_FAB2RAM_D1_I2, Tile_X9Y3_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_F (.I0(Tile_X9Y3_FAB2RAM_D1_I0), .I1(Tile_X9Y3_FAB2RAM_D1_I1), .I2(Tile_X9Y3_FAB2RAM_D1_I2), .I3(Tile_X9Y3_FAB2RAM_D1_I3));

wire Tile_X9Y3_FAB2RAM_D2_I0, Tile_X9Y3_FAB2RAM_D2_I1, Tile_X9Y3_FAB2RAM_D2_I2, Tile_X9Y3_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_G (.I0(Tile_X9Y3_FAB2RAM_D2_I0), .I1(Tile_X9Y3_FAB2RAM_D2_I1), .I2(Tile_X9Y3_FAB2RAM_D2_I2), .I3(Tile_X9Y3_FAB2RAM_D2_I3));

wire Tile_X9Y3_FAB2RAM_D3_I0, Tile_X9Y3_FAB2RAM_D3_I1, Tile_X9Y3_FAB2RAM_D3_I2, Tile_X9Y3_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_H (.I0(Tile_X9Y3_FAB2RAM_D3_I0), .I1(Tile_X9Y3_FAB2RAM_D3_I1), .I2(Tile_X9Y3_FAB2RAM_D3_I2), .I3(Tile_X9Y3_FAB2RAM_D3_I3));

wire Tile_X9Y3_FAB2RAM_A0_I0, Tile_X9Y3_FAB2RAM_A0_I1, Tile_X9Y3_FAB2RAM_A0_I2, Tile_X9Y3_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_I (.I0(Tile_X9Y3_FAB2RAM_A0_I0), .I1(Tile_X9Y3_FAB2RAM_A0_I1), .I2(Tile_X9Y3_FAB2RAM_A0_I2), .I3(Tile_X9Y3_FAB2RAM_A0_I3));

wire Tile_X9Y3_FAB2RAM_A1_I0, Tile_X9Y3_FAB2RAM_A1_I1, Tile_X9Y3_FAB2RAM_A1_I2, Tile_X9Y3_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_J (.I0(Tile_X9Y3_FAB2RAM_A1_I0), .I1(Tile_X9Y3_FAB2RAM_A1_I1), .I2(Tile_X9Y3_FAB2RAM_A1_I2), .I3(Tile_X9Y3_FAB2RAM_A1_I3));

wire Tile_X9Y3_FAB2RAM_C_I0, Tile_X9Y3_FAB2RAM_C_I1, Tile_X9Y3_FAB2RAM_C_I2, Tile_X9Y3_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y3_K (.I0(Tile_X9Y3_FAB2RAM_C_I0), .I1(Tile_X9Y3_FAB2RAM_C_I1), .I2(Tile_X9Y3_FAB2RAM_C_I2), .I3(Tile_X9Y3_FAB2RAM_C_I3));

wire Tile_X0Y4_A_I, Tile_X0Y4_A_T, Tile_X0Y4_A_O, Tile_X0Y4_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y4_A (.O(Tile_X0Y4_A_O), .Q(Tile_X0Y4_A_Q), .I(Tile_X0Y4_A_I));

wire Tile_X0Y4_B_I, Tile_X0Y4_B_T, Tile_X0Y4_B_O, Tile_X0Y4_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y4_B (.O(Tile_X0Y4_B_O), .Q(Tile_X0Y4_B_Q), .I(Tile_X0Y4_B_I));

wire Tile_X9Y4_RAM2FAB_D0_O0, Tile_X9Y4_RAM2FAB_D0_O1, Tile_X9Y4_RAM2FAB_D0_O2, Tile_X9Y4_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y4_A (.O0(Tile_X9Y4_RAM2FAB_D0_O0), .O1(Tile_X9Y4_RAM2FAB_D0_O1), .O2(Tile_X9Y4_RAM2FAB_D0_O2), .O3(Tile_X9Y4_RAM2FAB_D0_O3));

wire Tile_X9Y4_RAM2FAB_D1_O0, Tile_X9Y4_RAM2FAB_D1_O1, Tile_X9Y4_RAM2FAB_D1_O2, Tile_X9Y4_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y4_B (.O0(Tile_X9Y4_RAM2FAB_D1_O0), .O1(Tile_X9Y4_RAM2FAB_D1_O1), .O2(Tile_X9Y4_RAM2FAB_D1_O2), .O3(Tile_X9Y4_RAM2FAB_D1_O3));

wire Tile_X9Y4_RAM2FAB_D2_O0, Tile_X9Y4_RAM2FAB_D2_O1, Tile_X9Y4_RAM2FAB_D2_O2, Tile_X9Y4_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y4_C (.O0(Tile_X9Y4_RAM2FAB_D2_O0), .O1(Tile_X9Y4_RAM2FAB_D2_O1), .O2(Tile_X9Y4_RAM2FAB_D2_O2), .O3(Tile_X9Y4_RAM2FAB_D2_O3));

wire Tile_X9Y4_RAM2FAB_D3_O0, Tile_X9Y4_RAM2FAB_D3_O1, Tile_X9Y4_RAM2FAB_D3_O2, Tile_X9Y4_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y4_D (.O0(Tile_X9Y4_RAM2FAB_D3_O0), .O1(Tile_X9Y4_RAM2FAB_D3_O1), .O2(Tile_X9Y4_RAM2FAB_D3_O2), .O3(Tile_X9Y4_RAM2FAB_D3_O3));

wire Tile_X9Y4_FAB2RAM_D0_I0, Tile_X9Y4_FAB2RAM_D0_I1, Tile_X9Y4_FAB2RAM_D0_I2, Tile_X9Y4_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_E (.I0(Tile_X9Y4_FAB2RAM_D0_I0), .I1(Tile_X9Y4_FAB2RAM_D0_I1), .I2(Tile_X9Y4_FAB2RAM_D0_I2), .I3(Tile_X9Y4_FAB2RAM_D0_I3));

wire Tile_X9Y4_FAB2RAM_D1_I0, Tile_X9Y4_FAB2RAM_D1_I1, Tile_X9Y4_FAB2RAM_D1_I2, Tile_X9Y4_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_F (.I0(Tile_X9Y4_FAB2RAM_D1_I0), .I1(Tile_X9Y4_FAB2RAM_D1_I1), .I2(Tile_X9Y4_FAB2RAM_D1_I2), .I3(Tile_X9Y4_FAB2RAM_D1_I3));

wire Tile_X9Y4_FAB2RAM_D2_I0, Tile_X9Y4_FAB2RAM_D2_I1, Tile_X9Y4_FAB2RAM_D2_I2, Tile_X9Y4_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_G (.I0(Tile_X9Y4_FAB2RAM_D2_I0), .I1(Tile_X9Y4_FAB2RAM_D2_I1), .I2(Tile_X9Y4_FAB2RAM_D2_I2), .I3(Tile_X9Y4_FAB2RAM_D2_I3));

wire Tile_X9Y4_FAB2RAM_D3_I0, Tile_X9Y4_FAB2RAM_D3_I1, Tile_X9Y4_FAB2RAM_D3_I2, Tile_X9Y4_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_H (.I0(Tile_X9Y4_FAB2RAM_D3_I0), .I1(Tile_X9Y4_FAB2RAM_D3_I1), .I2(Tile_X9Y4_FAB2RAM_D3_I2), .I3(Tile_X9Y4_FAB2RAM_D3_I3));

wire Tile_X9Y4_FAB2RAM_A0_I0, Tile_X9Y4_FAB2RAM_A0_I1, Tile_X9Y4_FAB2RAM_A0_I2, Tile_X9Y4_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_I (.I0(Tile_X9Y4_FAB2RAM_A0_I0), .I1(Tile_X9Y4_FAB2RAM_A0_I1), .I2(Tile_X9Y4_FAB2RAM_A0_I2), .I3(Tile_X9Y4_FAB2RAM_A0_I3));

wire Tile_X9Y4_FAB2RAM_A1_I0, Tile_X9Y4_FAB2RAM_A1_I1, Tile_X9Y4_FAB2RAM_A1_I2, Tile_X9Y4_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_J (.I0(Tile_X9Y4_FAB2RAM_A1_I0), .I1(Tile_X9Y4_FAB2RAM_A1_I1), .I2(Tile_X9Y4_FAB2RAM_A1_I2), .I3(Tile_X9Y4_FAB2RAM_A1_I3));

wire Tile_X9Y4_FAB2RAM_C_I0, Tile_X9Y4_FAB2RAM_C_I1, Tile_X9Y4_FAB2RAM_C_I2, Tile_X9Y4_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y4_K (.I0(Tile_X9Y4_FAB2RAM_C_I0), .I1(Tile_X9Y4_FAB2RAM_C_I1), .I2(Tile_X9Y4_FAB2RAM_C_I2), .I3(Tile_X9Y4_FAB2RAM_C_I3));

wire Tile_X0Y5_A_I, Tile_X0Y5_A_T, Tile_X0Y5_A_O, Tile_X0Y5_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y5_A (.O(Tile_X0Y5_A_O), .Q(Tile_X0Y5_A_Q), .I(Tile_X0Y5_A_I));

wire Tile_X0Y5_B_I, Tile_X0Y5_B_T, Tile_X0Y5_B_O, Tile_X0Y5_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y5_B (.O(Tile_X0Y5_B_O), .Q(Tile_X0Y5_B_Q), .I(Tile_X0Y5_B_I));

wire Tile_X9Y5_RAM2FAB_D0_O0, Tile_X9Y5_RAM2FAB_D0_O1, Tile_X9Y5_RAM2FAB_D0_O2, Tile_X9Y5_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y5_A (.O0(Tile_X9Y5_RAM2FAB_D0_O0), .O1(Tile_X9Y5_RAM2FAB_D0_O1), .O2(Tile_X9Y5_RAM2FAB_D0_O2), .O3(Tile_X9Y5_RAM2FAB_D0_O3));

wire Tile_X9Y5_RAM2FAB_D1_O0, Tile_X9Y5_RAM2FAB_D1_O1, Tile_X9Y5_RAM2FAB_D1_O2, Tile_X9Y5_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y5_B (.O0(Tile_X9Y5_RAM2FAB_D1_O0), .O1(Tile_X9Y5_RAM2FAB_D1_O1), .O2(Tile_X9Y5_RAM2FAB_D1_O2), .O3(Tile_X9Y5_RAM2FAB_D1_O3));

wire Tile_X9Y5_RAM2FAB_D2_O0, Tile_X9Y5_RAM2FAB_D2_O1, Tile_X9Y5_RAM2FAB_D2_O2, Tile_X9Y5_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y5_C (.O0(Tile_X9Y5_RAM2FAB_D2_O0), .O1(Tile_X9Y5_RAM2FAB_D2_O1), .O2(Tile_X9Y5_RAM2FAB_D2_O2), .O3(Tile_X9Y5_RAM2FAB_D2_O3));

wire Tile_X9Y5_RAM2FAB_D3_O0, Tile_X9Y5_RAM2FAB_D3_O1, Tile_X9Y5_RAM2FAB_D3_O2, Tile_X9Y5_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y5_D (.O0(Tile_X9Y5_RAM2FAB_D3_O0), .O1(Tile_X9Y5_RAM2FAB_D3_O1), .O2(Tile_X9Y5_RAM2FAB_D3_O2), .O3(Tile_X9Y5_RAM2FAB_D3_O3));

wire Tile_X9Y5_FAB2RAM_D0_I0, Tile_X9Y5_FAB2RAM_D0_I1, Tile_X9Y5_FAB2RAM_D0_I2, Tile_X9Y5_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_E (.I0(Tile_X9Y5_FAB2RAM_D0_I0), .I1(Tile_X9Y5_FAB2RAM_D0_I1), .I2(Tile_X9Y5_FAB2RAM_D0_I2), .I3(Tile_X9Y5_FAB2RAM_D0_I3));

wire Tile_X9Y5_FAB2RAM_D1_I0, Tile_X9Y5_FAB2RAM_D1_I1, Tile_X9Y5_FAB2RAM_D1_I2, Tile_X9Y5_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_F (.I0(Tile_X9Y5_FAB2RAM_D1_I0), .I1(Tile_X9Y5_FAB2RAM_D1_I1), .I2(Tile_X9Y5_FAB2RAM_D1_I2), .I3(Tile_X9Y5_FAB2RAM_D1_I3));

wire Tile_X9Y5_FAB2RAM_D2_I0, Tile_X9Y5_FAB2RAM_D2_I1, Tile_X9Y5_FAB2RAM_D2_I2, Tile_X9Y5_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_G (.I0(Tile_X9Y5_FAB2RAM_D2_I0), .I1(Tile_X9Y5_FAB2RAM_D2_I1), .I2(Tile_X9Y5_FAB2RAM_D2_I2), .I3(Tile_X9Y5_FAB2RAM_D2_I3));

wire Tile_X9Y5_FAB2RAM_D3_I0, Tile_X9Y5_FAB2RAM_D3_I1, Tile_X9Y5_FAB2RAM_D3_I2, Tile_X9Y5_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_H (.I0(Tile_X9Y5_FAB2RAM_D3_I0), .I1(Tile_X9Y5_FAB2RAM_D3_I1), .I2(Tile_X9Y5_FAB2RAM_D3_I2), .I3(Tile_X9Y5_FAB2RAM_D3_I3));

wire Tile_X9Y5_FAB2RAM_A0_I0, Tile_X9Y5_FAB2RAM_A0_I1, Tile_X9Y5_FAB2RAM_A0_I2, Tile_X9Y5_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_I (.I0(Tile_X9Y5_FAB2RAM_A0_I0), .I1(Tile_X9Y5_FAB2RAM_A0_I1), .I2(Tile_X9Y5_FAB2RAM_A0_I2), .I3(Tile_X9Y5_FAB2RAM_A0_I3));

wire Tile_X9Y5_FAB2RAM_A1_I0, Tile_X9Y5_FAB2RAM_A1_I1, Tile_X9Y5_FAB2RAM_A1_I2, Tile_X9Y5_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_J (.I0(Tile_X9Y5_FAB2RAM_A1_I0), .I1(Tile_X9Y5_FAB2RAM_A1_I1), .I2(Tile_X9Y5_FAB2RAM_A1_I2), .I3(Tile_X9Y5_FAB2RAM_A1_I3));

wire Tile_X9Y5_FAB2RAM_C_I0, Tile_X9Y5_FAB2RAM_C_I1, Tile_X9Y5_FAB2RAM_C_I2, Tile_X9Y5_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y5_K (.I0(Tile_X9Y5_FAB2RAM_C_I0), .I1(Tile_X9Y5_FAB2RAM_C_I1), .I2(Tile_X9Y5_FAB2RAM_C_I2), .I3(Tile_X9Y5_FAB2RAM_C_I3));

wire Tile_X0Y6_A_I, Tile_X0Y6_A_T, Tile_X0Y6_A_O, Tile_X0Y6_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y6_A (.O(Tile_X0Y6_A_O), .Q(Tile_X0Y6_A_Q), .I(Tile_X0Y6_A_I));

wire Tile_X0Y6_B_I, Tile_X0Y6_B_T, Tile_X0Y6_B_O, Tile_X0Y6_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y6_B (.O(Tile_X0Y6_B_O), .Q(Tile_X0Y6_B_Q), .I(Tile_X0Y6_B_I));

wire Tile_X9Y6_RAM2FAB_D0_O0, Tile_X9Y6_RAM2FAB_D0_O1, Tile_X9Y6_RAM2FAB_D0_O2, Tile_X9Y6_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y6_A (.O0(Tile_X9Y6_RAM2FAB_D0_O0), .O1(Tile_X9Y6_RAM2FAB_D0_O1), .O2(Tile_X9Y6_RAM2FAB_D0_O2), .O3(Tile_X9Y6_RAM2FAB_D0_O3));

wire Tile_X9Y6_RAM2FAB_D1_O0, Tile_X9Y6_RAM2FAB_D1_O1, Tile_X9Y6_RAM2FAB_D1_O2, Tile_X9Y6_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y6_B (.O0(Tile_X9Y6_RAM2FAB_D1_O0), .O1(Tile_X9Y6_RAM2FAB_D1_O1), .O2(Tile_X9Y6_RAM2FAB_D1_O2), .O3(Tile_X9Y6_RAM2FAB_D1_O3));

wire Tile_X9Y6_RAM2FAB_D2_O0, Tile_X9Y6_RAM2FAB_D2_O1, Tile_X9Y6_RAM2FAB_D2_O2, Tile_X9Y6_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y6_C (.O0(Tile_X9Y6_RAM2FAB_D2_O0), .O1(Tile_X9Y6_RAM2FAB_D2_O1), .O2(Tile_X9Y6_RAM2FAB_D2_O2), .O3(Tile_X9Y6_RAM2FAB_D2_O3));

wire Tile_X9Y6_RAM2FAB_D3_O0, Tile_X9Y6_RAM2FAB_D3_O1, Tile_X9Y6_RAM2FAB_D3_O2, Tile_X9Y6_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y6_D (.O0(Tile_X9Y6_RAM2FAB_D3_O0), .O1(Tile_X9Y6_RAM2FAB_D3_O1), .O2(Tile_X9Y6_RAM2FAB_D3_O2), .O3(Tile_X9Y6_RAM2FAB_D3_O3));

wire Tile_X9Y6_FAB2RAM_D0_I0, Tile_X9Y6_FAB2RAM_D0_I1, Tile_X9Y6_FAB2RAM_D0_I2, Tile_X9Y6_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_E (.I0(Tile_X9Y6_FAB2RAM_D0_I0), .I1(Tile_X9Y6_FAB2RAM_D0_I1), .I2(Tile_X9Y6_FAB2RAM_D0_I2), .I3(Tile_X9Y6_FAB2RAM_D0_I3));

wire Tile_X9Y6_FAB2RAM_D1_I0, Tile_X9Y6_FAB2RAM_D1_I1, Tile_X9Y6_FAB2RAM_D1_I2, Tile_X9Y6_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_F (.I0(Tile_X9Y6_FAB2RAM_D1_I0), .I1(Tile_X9Y6_FAB2RAM_D1_I1), .I2(Tile_X9Y6_FAB2RAM_D1_I2), .I3(Tile_X9Y6_FAB2RAM_D1_I3));

wire Tile_X9Y6_FAB2RAM_D2_I0, Tile_X9Y6_FAB2RAM_D2_I1, Tile_X9Y6_FAB2RAM_D2_I2, Tile_X9Y6_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_G (.I0(Tile_X9Y6_FAB2RAM_D2_I0), .I1(Tile_X9Y6_FAB2RAM_D2_I1), .I2(Tile_X9Y6_FAB2RAM_D2_I2), .I3(Tile_X9Y6_FAB2RAM_D2_I3));

wire Tile_X9Y6_FAB2RAM_D3_I0, Tile_X9Y6_FAB2RAM_D3_I1, Tile_X9Y6_FAB2RAM_D3_I2, Tile_X9Y6_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_H (.I0(Tile_X9Y6_FAB2RAM_D3_I0), .I1(Tile_X9Y6_FAB2RAM_D3_I1), .I2(Tile_X9Y6_FAB2RAM_D3_I2), .I3(Tile_X9Y6_FAB2RAM_D3_I3));

wire Tile_X9Y6_FAB2RAM_A0_I0, Tile_X9Y6_FAB2RAM_A0_I1, Tile_X9Y6_FAB2RAM_A0_I2, Tile_X9Y6_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_I (.I0(Tile_X9Y6_FAB2RAM_A0_I0), .I1(Tile_X9Y6_FAB2RAM_A0_I1), .I2(Tile_X9Y6_FAB2RAM_A0_I2), .I3(Tile_X9Y6_FAB2RAM_A0_I3));

wire Tile_X9Y6_FAB2RAM_A1_I0, Tile_X9Y6_FAB2RAM_A1_I1, Tile_X9Y6_FAB2RAM_A1_I2, Tile_X9Y6_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_J (.I0(Tile_X9Y6_FAB2RAM_A1_I0), .I1(Tile_X9Y6_FAB2RAM_A1_I1), .I2(Tile_X9Y6_FAB2RAM_A1_I2), .I3(Tile_X9Y6_FAB2RAM_A1_I3));

wire Tile_X9Y6_FAB2RAM_C_I0, Tile_X9Y6_FAB2RAM_C_I1, Tile_X9Y6_FAB2RAM_C_I2, Tile_X9Y6_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y6_K (.I0(Tile_X9Y6_FAB2RAM_C_I0), .I1(Tile_X9Y6_FAB2RAM_C_I1), .I2(Tile_X9Y6_FAB2RAM_C_I2), .I3(Tile_X9Y6_FAB2RAM_C_I3));

wire Tile_X0Y7_A_I, Tile_X0Y7_A_T, Tile_X0Y7_A_O, Tile_X0Y7_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y7_A (.O(Tile_X0Y7_A_O), .Q(Tile_X0Y7_A_Q), .I(Tile_X0Y7_A_I));

wire Tile_X0Y7_B_I, Tile_X0Y7_B_T, Tile_X0Y7_B_O, Tile_X0Y7_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y7_B (.O(Tile_X0Y7_B_O), .Q(Tile_X0Y7_B_Q), .I(Tile_X0Y7_B_I));

wire Tile_X9Y7_RAM2FAB_D0_O0, Tile_X9Y7_RAM2FAB_D0_O1, Tile_X9Y7_RAM2FAB_D0_O2, Tile_X9Y7_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y7_A (.O0(Tile_X9Y7_RAM2FAB_D0_O0), .O1(Tile_X9Y7_RAM2FAB_D0_O1), .O2(Tile_X9Y7_RAM2FAB_D0_O2), .O3(Tile_X9Y7_RAM2FAB_D0_O3));

wire Tile_X9Y7_RAM2FAB_D1_O0, Tile_X9Y7_RAM2FAB_D1_O1, Tile_X9Y7_RAM2FAB_D1_O2, Tile_X9Y7_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y7_B (.O0(Tile_X9Y7_RAM2FAB_D1_O0), .O1(Tile_X9Y7_RAM2FAB_D1_O1), .O2(Tile_X9Y7_RAM2FAB_D1_O2), .O3(Tile_X9Y7_RAM2FAB_D1_O3));

wire Tile_X9Y7_RAM2FAB_D2_O0, Tile_X9Y7_RAM2FAB_D2_O1, Tile_X9Y7_RAM2FAB_D2_O2, Tile_X9Y7_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y7_C (.O0(Tile_X9Y7_RAM2FAB_D2_O0), .O1(Tile_X9Y7_RAM2FAB_D2_O1), .O2(Tile_X9Y7_RAM2FAB_D2_O2), .O3(Tile_X9Y7_RAM2FAB_D2_O3));

wire Tile_X9Y7_RAM2FAB_D3_O0, Tile_X9Y7_RAM2FAB_D3_O1, Tile_X9Y7_RAM2FAB_D3_O2, Tile_X9Y7_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y7_D (.O0(Tile_X9Y7_RAM2FAB_D3_O0), .O1(Tile_X9Y7_RAM2FAB_D3_O1), .O2(Tile_X9Y7_RAM2FAB_D3_O2), .O3(Tile_X9Y7_RAM2FAB_D3_O3));

wire Tile_X9Y7_FAB2RAM_D0_I0, Tile_X9Y7_FAB2RAM_D0_I1, Tile_X9Y7_FAB2RAM_D0_I2, Tile_X9Y7_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_E (.I0(Tile_X9Y7_FAB2RAM_D0_I0), .I1(Tile_X9Y7_FAB2RAM_D0_I1), .I2(Tile_X9Y7_FAB2RAM_D0_I2), .I3(Tile_X9Y7_FAB2RAM_D0_I3));

wire Tile_X9Y7_FAB2RAM_D1_I0, Tile_X9Y7_FAB2RAM_D1_I1, Tile_X9Y7_FAB2RAM_D1_I2, Tile_X9Y7_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_F (.I0(Tile_X9Y7_FAB2RAM_D1_I0), .I1(Tile_X9Y7_FAB2RAM_D1_I1), .I2(Tile_X9Y7_FAB2RAM_D1_I2), .I3(Tile_X9Y7_FAB2RAM_D1_I3));

wire Tile_X9Y7_FAB2RAM_D2_I0, Tile_X9Y7_FAB2RAM_D2_I1, Tile_X9Y7_FAB2RAM_D2_I2, Tile_X9Y7_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_G (.I0(Tile_X9Y7_FAB2RAM_D2_I0), .I1(Tile_X9Y7_FAB2RAM_D2_I1), .I2(Tile_X9Y7_FAB2RAM_D2_I2), .I3(Tile_X9Y7_FAB2RAM_D2_I3));

wire Tile_X9Y7_FAB2RAM_D3_I0, Tile_X9Y7_FAB2RAM_D3_I1, Tile_X9Y7_FAB2RAM_D3_I2, Tile_X9Y7_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_H (.I0(Tile_X9Y7_FAB2RAM_D3_I0), .I1(Tile_X9Y7_FAB2RAM_D3_I1), .I2(Tile_X9Y7_FAB2RAM_D3_I2), .I3(Tile_X9Y7_FAB2RAM_D3_I3));

wire Tile_X9Y7_FAB2RAM_A0_I0, Tile_X9Y7_FAB2RAM_A0_I1, Tile_X9Y7_FAB2RAM_A0_I2, Tile_X9Y7_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_I (.I0(Tile_X9Y7_FAB2RAM_A0_I0), .I1(Tile_X9Y7_FAB2RAM_A0_I1), .I2(Tile_X9Y7_FAB2RAM_A0_I2), .I3(Tile_X9Y7_FAB2RAM_A0_I3));

wire Tile_X9Y7_FAB2RAM_A1_I0, Tile_X9Y7_FAB2RAM_A1_I1, Tile_X9Y7_FAB2RAM_A1_I2, Tile_X9Y7_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_J (.I0(Tile_X9Y7_FAB2RAM_A1_I0), .I1(Tile_X9Y7_FAB2RAM_A1_I1), .I2(Tile_X9Y7_FAB2RAM_A1_I2), .I3(Tile_X9Y7_FAB2RAM_A1_I3));

wire Tile_X9Y7_FAB2RAM_C_I0, Tile_X9Y7_FAB2RAM_C_I1, Tile_X9Y7_FAB2RAM_C_I2, Tile_X9Y7_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y7_K (.I0(Tile_X9Y7_FAB2RAM_C_I0), .I1(Tile_X9Y7_FAB2RAM_C_I1), .I2(Tile_X9Y7_FAB2RAM_C_I2), .I3(Tile_X9Y7_FAB2RAM_C_I3));

wire Tile_X0Y8_A_I, Tile_X0Y8_A_T, Tile_X0Y8_A_O, Tile_X0Y8_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y8_A (.O(Tile_X0Y8_A_O), .Q(Tile_X0Y8_A_Q), .I(Tile_X0Y8_A_I));

wire Tile_X0Y8_B_I, Tile_X0Y8_B_T, Tile_X0Y8_B_O, Tile_X0Y8_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y8_B (.O(Tile_X0Y8_B_O), .Q(Tile_X0Y8_B_Q), .I(Tile_X0Y8_B_I));

wire Tile_X9Y8_RAM2FAB_D0_O0, Tile_X9Y8_RAM2FAB_D0_O1, Tile_X9Y8_RAM2FAB_D0_O2, Tile_X9Y8_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y8_A (.O0(Tile_X9Y8_RAM2FAB_D0_O0), .O1(Tile_X9Y8_RAM2FAB_D0_O1), .O2(Tile_X9Y8_RAM2FAB_D0_O2), .O3(Tile_X9Y8_RAM2FAB_D0_O3));

wire Tile_X9Y8_RAM2FAB_D1_O0, Tile_X9Y8_RAM2FAB_D1_O1, Tile_X9Y8_RAM2FAB_D1_O2, Tile_X9Y8_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y8_B (.O0(Tile_X9Y8_RAM2FAB_D1_O0), .O1(Tile_X9Y8_RAM2FAB_D1_O1), .O2(Tile_X9Y8_RAM2FAB_D1_O2), .O3(Tile_X9Y8_RAM2FAB_D1_O3));

wire Tile_X9Y8_RAM2FAB_D2_O0, Tile_X9Y8_RAM2FAB_D2_O1, Tile_X9Y8_RAM2FAB_D2_O2, Tile_X9Y8_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y8_C (.O0(Tile_X9Y8_RAM2FAB_D2_O0), .O1(Tile_X9Y8_RAM2FAB_D2_O1), .O2(Tile_X9Y8_RAM2FAB_D2_O2), .O3(Tile_X9Y8_RAM2FAB_D2_O3));

wire Tile_X9Y8_RAM2FAB_D3_O0, Tile_X9Y8_RAM2FAB_D3_O1, Tile_X9Y8_RAM2FAB_D3_O2, Tile_X9Y8_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y8_D (.O0(Tile_X9Y8_RAM2FAB_D3_O0), .O1(Tile_X9Y8_RAM2FAB_D3_O1), .O2(Tile_X9Y8_RAM2FAB_D3_O2), .O3(Tile_X9Y8_RAM2FAB_D3_O3));

wire Tile_X9Y8_FAB2RAM_D0_I0, Tile_X9Y8_FAB2RAM_D0_I1, Tile_X9Y8_FAB2RAM_D0_I2, Tile_X9Y8_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_E (.I0(Tile_X9Y8_FAB2RAM_D0_I0), .I1(Tile_X9Y8_FAB2RAM_D0_I1), .I2(Tile_X9Y8_FAB2RAM_D0_I2), .I3(Tile_X9Y8_FAB2RAM_D0_I3));

wire Tile_X9Y8_FAB2RAM_D1_I0, Tile_X9Y8_FAB2RAM_D1_I1, Tile_X9Y8_FAB2RAM_D1_I2, Tile_X9Y8_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_F (.I0(Tile_X9Y8_FAB2RAM_D1_I0), .I1(Tile_X9Y8_FAB2RAM_D1_I1), .I2(Tile_X9Y8_FAB2RAM_D1_I2), .I3(Tile_X9Y8_FAB2RAM_D1_I3));

wire Tile_X9Y8_FAB2RAM_D2_I0, Tile_X9Y8_FAB2RAM_D2_I1, Tile_X9Y8_FAB2RAM_D2_I2, Tile_X9Y8_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_G (.I0(Tile_X9Y8_FAB2RAM_D2_I0), .I1(Tile_X9Y8_FAB2RAM_D2_I1), .I2(Tile_X9Y8_FAB2RAM_D2_I2), .I3(Tile_X9Y8_FAB2RAM_D2_I3));

wire Tile_X9Y8_FAB2RAM_D3_I0, Tile_X9Y8_FAB2RAM_D3_I1, Tile_X9Y8_FAB2RAM_D3_I2, Tile_X9Y8_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_H (.I0(Tile_X9Y8_FAB2RAM_D3_I0), .I1(Tile_X9Y8_FAB2RAM_D3_I1), .I2(Tile_X9Y8_FAB2RAM_D3_I2), .I3(Tile_X9Y8_FAB2RAM_D3_I3));

wire Tile_X9Y8_FAB2RAM_A0_I0, Tile_X9Y8_FAB2RAM_A0_I1, Tile_X9Y8_FAB2RAM_A0_I2, Tile_X9Y8_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_I (.I0(Tile_X9Y8_FAB2RAM_A0_I0), .I1(Tile_X9Y8_FAB2RAM_A0_I1), .I2(Tile_X9Y8_FAB2RAM_A0_I2), .I3(Tile_X9Y8_FAB2RAM_A0_I3));

wire Tile_X9Y8_FAB2RAM_A1_I0, Tile_X9Y8_FAB2RAM_A1_I1, Tile_X9Y8_FAB2RAM_A1_I2, Tile_X9Y8_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_J (.I0(Tile_X9Y8_FAB2RAM_A1_I0), .I1(Tile_X9Y8_FAB2RAM_A1_I1), .I2(Tile_X9Y8_FAB2RAM_A1_I2), .I3(Tile_X9Y8_FAB2RAM_A1_I3));

wire Tile_X9Y8_FAB2RAM_C_I0, Tile_X9Y8_FAB2RAM_C_I1, Tile_X9Y8_FAB2RAM_C_I2, Tile_X9Y8_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y8_K (.I0(Tile_X9Y8_FAB2RAM_C_I0), .I1(Tile_X9Y8_FAB2RAM_C_I1), .I2(Tile_X9Y8_FAB2RAM_C_I2), .I3(Tile_X9Y8_FAB2RAM_C_I3));

wire Tile_X0Y9_A_I, Tile_X0Y9_A_T, Tile_X0Y9_A_O, Tile_X0Y9_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y9_A (.O(Tile_X0Y9_A_O), .Q(Tile_X0Y9_A_Q), .I(Tile_X0Y9_A_I));

wire Tile_X0Y9_B_I, Tile_X0Y9_B_T, Tile_X0Y9_B_O, Tile_X0Y9_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y9_B (.O(Tile_X0Y9_B_O), .Q(Tile_X0Y9_B_Q), .I(Tile_X0Y9_B_I));

wire Tile_X9Y9_RAM2FAB_D0_O0, Tile_X9Y9_RAM2FAB_D0_O1, Tile_X9Y9_RAM2FAB_D0_O2, Tile_X9Y9_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y9_A (.O0(Tile_X9Y9_RAM2FAB_D0_O0), .O1(Tile_X9Y9_RAM2FAB_D0_O1), .O2(Tile_X9Y9_RAM2FAB_D0_O2), .O3(Tile_X9Y9_RAM2FAB_D0_O3));

wire Tile_X9Y9_RAM2FAB_D1_O0, Tile_X9Y9_RAM2FAB_D1_O1, Tile_X9Y9_RAM2FAB_D1_O2, Tile_X9Y9_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y9_B (.O0(Tile_X9Y9_RAM2FAB_D1_O0), .O1(Tile_X9Y9_RAM2FAB_D1_O1), .O2(Tile_X9Y9_RAM2FAB_D1_O2), .O3(Tile_X9Y9_RAM2FAB_D1_O3));

wire Tile_X9Y9_RAM2FAB_D2_O0, Tile_X9Y9_RAM2FAB_D2_O1, Tile_X9Y9_RAM2FAB_D2_O2, Tile_X9Y9_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y9_C (.O0(Tile_X9Y9_RAM2FAB_D2_O0), .O1(Tile_X9Y9_RAM2FAB_D2_O1), .O2(Tile_X9Y9_RAM2FAB_D2_O2), .O3(Tile_X9Y9_RAM2FAB_D2_O3));

wire Tile_X9Y9_RAM2FAB_D3_O0, Tile_X9Y9_RAM2FAB_D3_O1, Tile_X9Y9_RAM2FAB_D3_O2, Tile_X9Y9_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y9_D (.O0(Tile_X9Y9_RAM2FAB_D3_O0), .O1(Tile_X9Y9_RAM2FAB_D3_O1), .O2(Tile_X9Y9_RAM2FAB_D3_O2), .O3(Tile_X9Y9_RAM2FAB_D3_O3));

wire Tile_X9Y9_FAB2RAM_D0_I0, Tile_X9Y9_FAB2RAM_D0_I1, Tile_X9Y9_FAB2RAM_D0_I2, Tile_X9Y9_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_E (.I0(Tile_X9Y9_FAB2RAM_D0_I0), .I1(Tile_X9Y9_FAB2RAM_D0_I1), .I2(Tile_X9Y9_FAB2RAM_D0_I2), .I3(Tile_X9Y9_FAB2RAM_D0_I3));

wire Tile_X9Y9_FAB2RAM_D1_I0, Tile_X9Y9_FAB2RAM_D1_I1, Tile_X9Y9_FAB2RAM_D1_I2, Tile_X9Y9_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_F (.I0(Tile_X9Y9_FAB2RAM_D1_I0), .I1(Tile_X9Y9_FAB2RAM_D1_I1), .I2(Tile_X9Y9_FAB2RAM_D1_I2), .I3(Tile_X9Y9_FAB2RAM_D1_I3));

wire Tile_X9Y9_FAB2RAM_D2_I0, Tile_X9Y9_FAB2RAM_D2_I1, Tile_X9Y9_FAB2RAM_D2_I2, Tile_X9Y9_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_G (.I0(Tile_X9Y9_FAB2RAM_D2_I0), .I1(Tile_X9Y9_FAB2RAM_D2_I1), .I2(Tile_X9Y9_FAB2RAM_D2_I2), .I3(Tile_X9Y9_FAB2RAM_D2_I3));

wire Tile_X9Y9_FAB2RAM_D3_I0, Tile_X9Y9_FAB2RAM_D3_I1, Tile_X9Y9_FAB2RAM_D3_I2, Tile_X9Y9_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_H (.I0(Tile_X9Y9_FAB2RAM_D3_I0), .I1(Tile_X9Y9_FAB2RAM_D3_I1), .I2(Tile_X9Y9_FAB2RAM_D3_I2), .I3(Tile_X9Y9_FAB2RAM_D3_I3));

wire Tile_X9Y9_FAB2RAM_A0_I0, Tile_X9Y9_FAB2RAM_A0_I1, Tile_X9Y9_FAB2RAM_A0_I2, Tile_X9Y9_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_I (.I0(Tile_X9Y9_FAB2RAM_A0_I0), .I1(Tile_X9Y9_FAB2RAM_A0_I1), .I2(Tile_X9Y9_FAB2RAM_A0_I2), .I3(Tile_X9Y9_FAB2RAM_A0_I3));

wire Tile_X9Y9_FAB2RAM_A1_I0, Tile_X9Y9_FAB2RAM_A1_I1, Tile_X9Y9_FAB2RAM_A1_I2, Tile_X9Y9_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_J (.I0(Tile_X9Y9_FAB2RAM_A1_I0), .I1(Tile_X9Y9_FAB2RAM_A1_I1), .I2(Tile_X9Y9_FAB2RAM_A1_I2), .I3(Tile_X9Y9_FAB2RAM_A1_I3));

wire Tile_X9Y9_FAB2RAM_C_I0, Tile_X9Y9_FAB2RAM_C_I1, Tile_X9Y9_FAB2RAM_C_I2, Tile_X9Y9_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y9_K (.I0(Tile_X9Y9_FAB2RAM_C_I0), .I1(Tile_X9Y9_FAB2RAM_C_I1), .I2(Tile_X9Y9_FAB2RAM_C_I2), .I3(Tile_X9Y9_FAB2RAM_C_I3));

wire Tile_X0Y10_A_I, Tile_X0Y10_A_T, Tile_X0Y10_A_O, Tile_X0Y10_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_A (.O(Tile_X0Y10_A_O), .Q(Tile_X0Y10_A_Q), .I(Tile_X0Y10_A_I));

wire Tile_X0Y10_B_I, Tile_X0Y10_B_T, Tile_X0Y10_B_O, Tile_X0Y10_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_B (.O(Tile_X0Y10_B_O), .Q(Tile_X0Y10_B_Q), .I(Tile_X0Y10_B_I));

wire Tile_X9Y10_RAM2FAB_D0_O0, Tile_X9Y10_RAM2FAB_D0_O1, Tile_X9Y10_RAM2FAB_D0_O2, Tile_X9Y10_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y10_A (.O0(Tile_X9Y10_RAM2FAB_D0_O0), .O1(Tile_X9Y10_RAM2FAB_D0_O1), .O2(Tile_X9Y10_RAM2FAB_D0_O2), .O3(Tile_X9Y10_RAM2FAB_D0_O3));

wire Tile_X9Y10_RAM2FAB_D1_O0, Tile_X9Y10_RAM2FAB_D1_O1, Tile_X9Y10_RAM2FAB_D1_O2, Tile_X9Y10_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y10_B (.O0(Tile_X9Y10_RAM2FAB_D1_O0), .O1(Tile_X9Y10_RAM2FAB_D1_O1), .O2(Tile_X9Y10_RAM2FAB_D1_O2), .O3(Tile_X9Y10_RAM2FAB_D1_O3));

wire Tile_X9Y10_RAM2FAB_D2_O0, Tile_X9Y10_RAM2FAB_D2_O1, Tile_X9Y10_RAM2FAB_D2_O2, Tile_X9Y10_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y10_C (.O0(Tile_X9Y10_RAM2FAB_D2_O0), .O1(Tile_X9Y10_RAM2FAB_D2_O1), .O2(Tile_X9Y10_RAM2FAB_D2_O2), .O3(Tile_X9Y10_RAM2FAB_D2_O3));

wire Tile_X9Y10_RAM2FAB_D3_O0, Tile_X9Y10_RAM2FAB_D3_O1, Tile_X9Y10_RAM2FAB_D3_O2, Tile_X9Y10_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y10_D (.O0(Tile_X9Y10_RAM2FAB_D3_O0), .O1(Tile_X9Y10_RAM2FAB_D3_O1), .O2(Tile_X9Y10_RAM2FAB_D3_O2), .O3(Tile_X9Y10_RAM2FAB_D3_O3));

wire Tile_X9Y10_FAB2RAM_D0_I0, Tile_X9Y10_FAB2RAM_D0_I1, Tile_X9Y10_FAB2RAM_D0_I2, Tile_X9Y10_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_E (.I0(Tile_X9Y10_FAB2RAM_D0_I0), .I1(Tile_X9Y10_FAB2RAM_D0_I1), .I2(Tile_X9Y10_FAB2RAM_D0_I2), .I3(Tile_X9Y10_FAB2RAM_D0_I3));

wire Tile_X9Y10_FAB2RAM_D1_I0, Tile_X9Y10_FAB2RAM_D1_I1, Tile_X9Y10_FAB2RAM_D1_I2, Tile_X9Y10_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_F (.I0(Tile_X9Y10_FAB2RAM_D1_I0), .I1(Tile_X9Y10_FAB2RAM_D1_I1), .I2(Tile_X9Y10_FAB2RAM_D1_I2), .I3(Tile_X9Y10_FAB2RAM_D1_I3));

wire Tile_X9Y10_FAB2RAM_D2_I0, Tile_X9Y10_FAB2RAM_D2_I1, Tile_X9Y10_FAB2RAM_D2_I2, Tile_X9Y10_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_G (.I0(Tile_X9Y10_FAB2RAM_D2_I0), .I1(Tile_X9Y10_FAB2RAM_D2_I1), .I2(Tile_X9Y10_FAB2RAM_D2_I2), .I3(Tile_X9Y10_FAB2RAM_D2_I3));

wire Tile_X9Y10_FAB2RAM_D3_I0, Tile_X9Y10_FAB2RAM_D3_I1, Tile_X9Y10_FAB2RAM_D3_I2, Tile_X9Y10_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_H (.I0(Tile_X9Y10_FAB2RAM_D3_I0), .I1(Tile_X9Y10_FAB2RAM_D3_I1), .I2(Tile_X9Y10_FAB2RAM_D3_I2), .I3(Tile_X9Y10_FAB2RAM_D3_I3));

wire Tile_X9Y10_FAB2RAM_A0_I0, Tile_X9Y10_FAB2RAM_A0_I1, Tile_X9Y10_FAB2RAM_A0_I2, Tile_X9Y10_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_I (.I0(Tile_X9Y10_FAB2RAM_A0_I0), .I1(Tile_X9Y10_FAB2RAM_A0_I1), .I2(Tile_X9Y10_FAB2RAM_A0_I2), .I3(Tile_X9Y10_FAB2RAM_A0_I3));

wire Tile_X9Y10_FAB2RAM_A1_I0, Tile_X9Y10_FAB2RAM_A1_I1, Tile_X9Y10_FAB2RAM_A1_I2, Tile_X9Y10_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_J (.I0(Tile_X9Y10_FAB2RAM_A1_I0), .I1(Tile_X9Y10_FAB2RAM_A1_I1), .I2(Tile_X9Y10_FAB2RAM_A1_I2), .I3(Tile_X9Y10_FAB2RAM_A1_I3));

wire Tile_X9Y10_FAB2RAM_C_I0, Tile_X9Y10_FAB2RAM_C_I1, Tile_X9Y10_FAB2RAM_C_I2, Tile_X9Y10_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y10_K (.I0(Tile_X9Y10_FAB2RAM_C_I0), .I1(Tile_X9Y10_FAB2RAM_C_I1), .I2(Tile_X9Y10_FAB2RAM_C_I2), .I3(Tile_X9Y10_FAB2RAM_C_I3));

wire Tile_X0Y11_A_I, Tile_X0Y11_A_T, Tile_X0Y11_A_O, Tile_X0Y11_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_A (.O(Tile_X0Y11_A_O), .Q(Tile_X0Y11_A_Q), .I(Tile_X0Y11_A_I));

wire Tile_X0Y11_B_I, Tile_X0Y11_B_T, Tile_X0Y11_B_O, Tile_X0Y11_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_B (.O(Tile_X0Y11_B_O), .Q(Tile_X0Y11_B_Q), .I(Tile_X0Y11_B_I));

wire Tile_X9Y11_RAM2FAB_D0_O0, Tile_X9Y11_RAM2FAB_D0_O1, Tile_X9Y11_RAM2FAB_D0_O2, Tile_X9Y11_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y11_A (.O0(Tile_X9Y11_RAM2FAB_D0_O0), .O1(Tile_X9Y11_RAM2FAB_D0_O1), .O2(Tile_X9Y11_RAM2FAB_D0_O2), .O3(Tile_X9Y11_RAM2FAB_D0_O3));

wire Tile_X9Y11_RAM2FAB_D1_O0, Tile_X9Y11_RAM2FAB_D1_O1, Tile_X9Y11_RAM2FAB_D1_O2, Tile_X9Y11_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y11_B (.O0(Tile_X9Y11_RAM2FAB_D1_O0), .O1(Tile_X9Y11_RAM2FAB_D1_O1), .O2(Tile_X9Y11_RAM2FAB_D1_O2), .O3(Tile_X9Y11_RAM2FAB_D1_O3));

wire Tile_X9Y11_RAM2FAB_D2_O0, Tile_X9Y11_RAM2FAB_D2_O1, Tile_X9Y11_RAM2FAB_D2_O2, Tile_X9Y11_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y11_C (.O0(Tile_X9Y11_RAM2FAB_D2_O0), .O1(Tile_X9Y11_RAM2FAB_D2_O1), .O2(Tile_X9Y11_RAM2FAB_D2_O2), .O3(Tile_X9Y11_RAM2FAB_D2_O3));

wire Tile_X9Y11_RAM2FAB_D3_O0, Tile_X9Y11_RAM2FAB_D3_O1, Tile_X9Y11_RAM2FAB_D3_O2, Tile_X9Y11_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y11_D (.O0(Tile_X9Y11_RAM2FAB_D3_O0), .O1(Tile_X9Y11_RAM2FAB_D3_O1), .O2(Tile_X9Y11_RAM2FAB_D3_O2), .O3(Tile_X9Y11_RAM2FAB_D3_O3));

wire Tile_X9Y11_FAB2RAM_D0_I0, Tile_X9Y11_FAB2RAM_D0_I1, Tile_X9Y11_FAB2RAM_D0_I2, Tile_X9Y11_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_E (.I0(Tile_X9Y11_FAB2RAM_D0_I0), .I1(Tile_X9Y11_FAB2RAM_D0_I1), .I2(Tile_X9Y11_FAB2RAM_D0_I2), .I3(Tile_X9Y11_FAB2RAM_D0_I3));

wire Tile_X9Y11_FAB2RAM_D1_I0, Tile_X9Y11_FAB2RAM_D1_I1, Tile_X9Y11_FAB2RAM_D1_I2, Tile_X9Y11_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_F (.I0(Tile_X9Y11_FAB2RAM_D1_I0), .I1(Tile_X9Y11_FAB2RAM_D1_I1), .I2(Tile_X9Y11_FAB2RAM_D1_I2), .I3(Tile_X9Y11_FAB2RAM_D1_I3));

wire Tile_X9Y11_FAB2RAM_D2_I0, Tile_X9Y11_FAB2RAM_D2_I1, Tile_X9Y11_FAB2RAM_D2_I2, Tile_X9Y11_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_G (.I0(Tile_X9Y11_FAB2RAM_D2_I0), .I1(Tile_X9Y11_FAB2RAM_D2_I1), .I2(Tile_X9Y11_FAB2RAM_D2_I2), .I3(Tile_X9Y11_FAB2RAM_D2_I3));

wire Tile_X9Y11_FAB2RAM_D3_I0, Tile_X9Y11_FAB2RAM_D3_I1, Tile_X9Y11_FAB2RAM_D3_I2, Tile_X9Y11_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_H (.I0(Tile_X9Y11_FAB2RAM_D3_I0), .I1(Tile_X9Y11_FAB2RAM_D3_I1), .I2(Tile_X9Y11_FAB2RAM_D3_I2), .I3(Tile_X9Y11_FAB2RAM_D3_I3));

wire Tile_X9Y11_FAB2RAM_A0_I0, Tile_X9Y11_FAB2RAM_A0_I1, Tile_X9Y11_FAB2RAM_A0_I2, Tile_X9Y11_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_I (.I0(Tile_X9Y11_FAB2RAM_A0_I0), .I1(Tile_X9Y11_FAB2RAM_A0_I1), .I2(Tile_X9Y11_FAB2RAM_A0_I2), .I3(Tile_X9Y11_FAB2RAM_A0_I3));

wire Tile_X9Y11_FAB2RAM_A1_I0, Tile_X9Y11_FAB2RAM_A1_I1, Tile_X9Y11_FAB2RAM_A1_I2, Tile_X9Y11_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_J (.I0(Tile_X9Y11_FAB2RAM_A1_I0), .I1(Tile_X9Y11_FAB2RAM_A1_I1), .I2(Tile_X9Y11_FAB2RAM_A1_I2), .I3(Tile_X9Y11_FAB2RAM_A1_I3));

wire Tile_X9Y11_FAB2RAM_C_I0, Tile_X9Y11_FAB2RAM_C_I1, Tile_X9Y11_FAB2RAM_C_I2, Tile_X9Y11_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y11_K (.I0(Tile_X9Y11_FAB2RAM_C_I0), .I1(Tile_X9Y11_FAB2RAM_C_I1), .I2(Tile_X9Y11_FAB2RAM_C_I2), .I3(Tile_X9Y11_FAB2RAM_C_I3));

wire Tile_X0Y12_A_I, Tile_X0Y12_A_T, Tile_X0Y12_A_O, Tile_X0Y12_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_A (.O(Tile_X0Y12_A_O), .Q(Tile_X0Y12_A_Q), .I(Tile_X0Y12_A_I));

wire Tile_X0Y12_B_I, Tile_X0Y12_B_T, Tile_X0Y12_B_O, Tile_X0Y12_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_B (.O(Tile_X0Y12_B_O), .Q(Tile_X0Y12_B_Q), .I(Tile_X0Y12_B_I));

wire Tile_X9Y12_RAM2FAB_D0_O0, Tile_X9Y12_RAM2FAB_D0_O1, Tile_X9Y12_RAM2FAB_D0_O2, Tile_X9Y12_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X9Y12_A (.O0(Tile_X9Y12_RAM2FAB_D0_O0), .O1(Tile_X9Y12_RAM2FAB_D0_O1), .O2(Tile_X9Y12_RAM2FAB_D0_O2), .O3(Tile_X9Y12_RAM2FAB_D0_O3));

wire Tile_X9Y12_RAM2FAB_D1_O0, Tile_X9Y12_RAM2FAB_D1_O1, Tile_X9Y12_RAM2FAB_D1_O2, Tile_X9Y12_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X9Y12_B (.O0(Tile_X9Y12_RAM2FAB_D1_O0), .O1(Tile_X9Y12_RAM2FAB_D1_O1), .O2(Tile_X9Y12_RAM2FAB_D1_O2), .O3(Tile_X9Y12_RAM2FAB_D1_O3));

wire Tile_X9Y12_RAM2FAB_D2_O0, Tile_X9Y12_RAM2FAB_D2_O1, Tile_X9Y12_RAM2FAB_D2_O2, Tile_X9Y12_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X9Y12_C (.O0(Tile_X9Y12_RAM2FAB_D2_O0), .O1(Tile_X9Y12_RAM2FAB_D2_O1), .O2(Tile_X9Y12_RAM2FAB_D2_O2), .O3(Tile_X9Y12_RAM2FAB_D2_O3));

wire Tile_X9Y12_RAM2FAB_D3_O0, Tile_X9Y12_RAM2FAB_D3_O1, Tile_X9Y12_RAM2FAB_D3_O2, Tile_X9Y12_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X9Y12_D (.O0(Tile_X9Y12_RAM2FAB_D3_O0), .O1(Tile_X9Y12_RAM2FAB_D3_O1), .O2(Tile_X9Y12_RAM2FAB_D3_O2), .O3(Tile_X9Y12_RAM2FAB_D3_O3));

wire Tile_X9Y12_FAB2RAM_D0_I0, Tile_X9Y12_FAB2RAM_D0_I1, Tile_X9Y12_FAB2RAM_D0_I2, Tile_X9Y12_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_E (.I0(Tile_X9Y12_FAB2RAM_D0_I0), .I1(Tile_X9Y12_FAB2RAM_D0_I1), .I2(Tile_X9Y12_FAB2RAM_D0_I2), .I3(Tile_X9Y12_FAB2RAM_D0_I3));

wire Tile_X9Y12_FAB2RAM_D1_I0, Tile_X9Y12_FAB2RAM_D1_I1, Tile_X9Y12_FAB2RAM_D1_I2, Tile_X9Y12_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_F (.I0(Tile_X9Y12_FAB2RAM_D1_I0), .I1(Tile_X9Y12_FAB2RAM_D1_I1), .I2(Tile_X9Y12_FAB2RAM_D1_I2), .I3(Tile_X9Y12_FAB2RAM_D1_I3));

wire Tile_X9Y12_FAB2RAM_D2_I0, Tile_X9Y12_FAB2RAM_D2_I1, Tile_X9Y12_FAB2RAM_D2_I2, Tile_X9Y12_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_G (.I0(Tile_X9Y12_FAB2RAM_D2_I0), .I1(Tile_X9Y12_FAB2RAM_D2_I1), .I2(Tile_X9Y12_FAB2RAM_D2_I2), .I3(Tile_X9Y12_FAB2RAM_D2_I3));

wire Tile_X9Y12_FAB2RAM_D3_I0, Tile_X9Y12_FAB2RAM_D3_I1, Tile_X9Y12_FAB2RAM_D3_I2, Tile_X9Y12_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_H (.I0(Tile_X9Y12_FAB2RAM_D3_I0), .I1(Tile_X9Y12_FAB2RAM_D3_I1), .I2(Tile_X9Y12_FAB2RAM_D3_I2), .I3(Tile_X9Y12_FAB2RAM_D3_I3));

wire Tile_X9Y12_FAB2RAM_A0_I0, Tile_X9Y12_FAB2RAM_A0_I1, Tile_X9Y12_FAB2RAM_A0_I2, Tile_X9Y12_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_I (.I0(Tile_X9Y12_FAB2RAM_A0_I0), .I1(Tile_X9Y12_FAB2RAM_A0_I1), .I2(Tile_X9Y12_FAB2RAM_A0_I2), .I3(Tile_X9Y12_FAB2RAM_A0_I3));

wire Tile_X9Y12_FAB2RAM_A1_I0, Tile_X9Y12_FAB2RAM_A1_I1, Tile_X9Y12_FAB2RAM_A1_I2, Tile_X9Y12_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_J (.I0(Tile_X9Y12_FAB2RAM_A1_I0), .I1(Tile_X9Y12_FAB2RAM_A1_I1), .I2(Tile_X9Y12_FAB2RAM_A1_I2), .I3(Tile_X9Y12_FAB2RAM_A1_I3));

wire Tile_X9Y12_FAB2RAM_C_I0, Tile_X9Y12_FAB2RAM_C_I1, Tile_X9Y12_FAB2RAM_C_I2, Tile_X9Y12_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X9Y12_K (.I0(Tile_X9Y12_FAB2RAM_C_I0), .I1(Tile_X9Y12_FAB2RAM_C_I1), .I2(Tile_X9Y12_FAB2RAM_C_I2), .I3(Tile_X9Y12_FAB2RAM_C_I3));

endmodule